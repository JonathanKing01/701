// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.0 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Mon May  6 09:14:11 2019
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [3:0] LEGUP_0 = 4'd0;
parameter [3:0] LEGUP_F_main_BB_entry_1 = 4'd1;
parameter [3:0] LEGUP_pipeline_wait_loop_2 = 4'd2;
parameter [3:0] LEGUP_F_main_BB_for_cond2_preheader_preheader_3 = 4'd3;
parameter [3:0] LEGUP_F_main_BB_for_cond2_preheader_preheader_4 = 4'd4;
parameter [3:0] LEGUP_F_main_BB_for_cond2_preheader_preheader_5 = 4'd5;
parameter [3:0] LEGUP_F_main_BB_for_cond2_preheader_preheader_6 = 4'd6;
parameter [3:0] LEGUP_F_main_BB_for_cond2_preheader_preheader_7 = 4'd7;
parameter [3:0] LEGUP_F_main_BB_for_cond2_preheader_8 = 4'd8;
parameter [3:0] LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9 = 4'd9;
parameter [3:0] LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10 = 4'd10;
parameter [3:0] LEGUP_F_main_BB_for_end9_11 = 4'd11;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [3:0] cur_state;
reg [3:0] next_state;
wire  fsm_stall;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_0;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_0_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_1;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_1_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_2_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_4_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_5_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_6_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_7;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_8_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_9;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_10;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_11;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_11_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_12;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_12_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_13;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_13_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_14;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_14_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_15;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_15_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_16;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_17;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_17_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_18;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_18_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_19;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_19_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_20;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_20_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_21;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_22_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_23;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_24;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_24_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_25;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_25_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_26;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_26_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_27;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_27_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_28;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_29;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_29_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_30;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_30_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_31;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_32;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_32_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_33;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_33_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_34;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_34_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_35;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_36;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_36_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_37;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_37_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_38;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_39;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_39_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_40;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_40_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_41;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_41_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_42;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_43;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_43_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_44;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_44_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_45;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_46;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_46_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_47;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_47_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_48;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_48_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_49;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_50;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_50_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_51;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_51_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_52;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_53;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_53_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_54;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_54_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_55;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_55_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_preheader_56;
reg [31:0] main_for_cond2_preheader_57;
reg [31:0] main_for_cond2_preheader_57_reg;
reg [31:0] main_for_cond2_preheader_58;
reg [31:0] main_for_cond2_preheader_58_reg;
reg [31:0] main_for_cond2_preheader_59;
reg [31:0] main_for_cond2_preheader_59_reg;
reg [31:0] main_for_cond2_preheader_60;
reg [31:0] main_for_cond2_preheader_60_reg;
reg [31:0] main_for_cond2_preheader_61;
reg [31:0] main_for_cond2_preheader_61_reg;
reg [31:0] main_for_cond2_preheader_62;
reg [31:0] main_for_cond2_preheader_62_reg;
reg [31:0] main_for_cond2_preheader_63;
reg [31:0] main_for_cond2_preheader_63_reg;
reg [31:0] main_for_cond2_preheader_64;
reg [31:0] main_for_cond2_preheader_64_reg;
reg [3:0] main_for_cond2_preheader_65;
reg [3:0] main_for_cond2_preheader_65_reg;
reg  main_for_cond2_preheader_exitcond1;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_for_cond2_preheader_crit_;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_for_cond2_preheader_crit__var0;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_for_cond2_preheader_crit__var1;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_for_cond2_preheader_crit__var2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_for_cond2_preheader_crit__var3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_for_cond2_preheader_crit__var4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_for_cond2_preheader_crit__var5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond2_preheader_for_cond2_preheader_crit__var6;
reg [4:0] main_for_cond2_preheader_for_cond2_preheader_crit__var7;
reg [4:0] main_for_cond2_preheader_for_cond2_preheader_crit__var7_reg;
reg [31:0] main_for_cond2_preheader_for_cond2_preheader_crit__var8;
reg [31:0] main_for_cond2_preheader_for_cond2_preheader_crit__var9;
reg [31:0] main_for_cond2_preheader_for_cond2_preheader_crit__var10;
reg [31:0] main_for_cond2_preheader_for_cond2_preheader_crit__var11;
reg [31:0] main_for_cond2_preheader_for_cond2_preheader_crit__var12;
reg [31:0] main_for_cond2_preheader_for_cond2_preheader_crit__var13;
reg [31:0] main_for_cond2_preheader_for_cond2_preheader_crit__var14;
reg [31:0] main_for_cond2_preheader_for_cond2_preheader_crit__var15;
reg [2:0] main_entry_DCT1_address_a;
reg  main_entry_DCT1_write_enable_a;
reg [31:0] main_entry_DCT1_in_a;
wire [31:0] main_entry_DCT1_out_a;
reg [2:0] main_entry_DCT1_address_b;
reg  main_entry_DCT1_write_enable_b;
reg [31:0] main_entry_DCT1_in_b;
wire [31:0] main_entry_DCT1_out_b;
reg [2:0] main_entry_DCT2_address_a;
reg  main_entry_DCT2_write_enable_a;
reg [31:0] main_entry_DCT2_in_a;
wire [31:0] main_entry_DCT2_out_a;
reg [2:0] main_entry_DCT2_address_b;
reg  main_entry_DCT2_write_enable_b;
reg [31:0] main_entry_DCT2_in_b;
wire [31:0] main_entry_DCT2_out_b;
reg [2:0] main_entry_DCT3_address_a;
reg  main_entry_DCT3_write_enable_a;
reg [31:0] main_entry_DCT3_in_a;
wire [31:0] main_entry_DCT3_out_a;
reg [2:0] main_entry_DCT3_address_b;
reg  main_entry_DCT3_write_enable_b;
reg [31:0] main_entry_DCT3_in_b;
wire [31:0] main_entry_DCT3_out_b;
reg [2:0] main_entry_DCT4_address_a;
reg  main_entry_DCT4_write_enable_a;
reg [31:0] main_entry_DCT4_in_a;
wire [31:0] main_entry_DCT4_out_a;
reg [2:0] main_entry_DCT4_address_b;
reg  main_entry_DCT4_write_enable_b;
reg [31:0] main_entry_DCT4_in_b;
wire [31:0] main_entry_DCT4_out_b;
reg [2:0] main_entry_DCT5_address_a;
reg  main_entry_DCT5_write_enable_a;
reg [31:0] main_entry_DCT5_in_a;
wire [31:0] main_entry_DCT5_out_a;
reg [2:0] main_entry_DCT5_address_b;
reg  main_entry_DCT5_write_enable_b;
reg [31:0] main_entry_DCT5_in_b;
wire [31:0] main_entry_DCT5_out_b;
reg [2:0] main_entry_DCT6_address_a;
reg  main_entry_DCT6_write_enable_a;
reg [31:0] main_entry_DCT6_in_a;
wire [31:0] main_entry_DCT6_out_a;
reg [2:0] main_entry_DCT6_address_b;
reg  main_entry_DCT6_write_enable_b;
reg [31:0] main_entry_DCT6_in_b;
wire [31:0] main_entry_DCT6_out_b;
reg [2:0] main_entry_DCT7_address_a;
reg  main_entry_DCT7_write_enable_a;
reg [31:0] main_entry_DCT7_in_a;
wire [31:0] main_entry_DCT7_out_a;
reg [2:0] main_entry_DCT7_address_b;
reg  main_entry_DCT7_write_enable_b;
reg [31:0] main_entry_DCT7_in_b;
wire [31:0] main_entry_DCT7_out_b;
reg [2:0] main_entry_DCT8_address_a;
reg  main_entry_DCT8_write_enable_a;
reg [31:0] main_entry_DCT8_in_a;
wire [31:0] main_entry_DCT8_out_a;
reg [2:0] main_entry_DCT8_address_b;
reg  main_entry_DCT8_write_enable_b;
reg [31:0] main_entry_DCT8_in_b;
wire [31:0] main_entry_DCT8_out_b;
reg  loop_valid_bit_0;
wire  loop_state_stall_0;
reg  loop_state_enable_0;
reg  loop_II_counter;
reg  loop_start;
reg  loop_activate_pipeline;
reg  loop_pipeline_exit_cond;
reg [31:0] loop_inductionVar_stage0;
reg  loop_active;
reg  loop_begin_pipeline;
reg  loop_epilogue;
reg  loop_pipeline_finish;
reg  loop_only_last_stage_enabled;
reg  loop_pipeline_finish_reg;



//   %DCT1 = alloca [7 x i32], align 4, !MSB !129, !LSB !130, !extendFrom !129
ram_dual_port main_entry_DCT1 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_DCT1_address_a ),
	.wren_a( main_entry_DCT1_write_enable_a ),
	.data_a( main_entry_DCT1_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_DCT1_out_a ),
	.address_b( main_entry_DCT1_address_b ),
	.wren_b( main_entry_DCT1_write_enable_b ),
	.data_b( main_entry_DCT1_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_DCT1_out_b )
);
defparam main_entry_DCT1.width_a = 32;
defparam main_entry_DCT1.widthad_a = 3;
defparam main_entry_DCT1.width_be_a = 4;
defparam main_entry_DCT1.numwords_a = 7;
defparam main_entry_DCT1.width_b = 32;
defparam main_entry_DCT1.widthad_b = 3;
defparam main_entry_DCT1.width_be_b = 4;
defparam main_entry_DCT1.numwords_b = 7;
defparam main_entry_DCT1.latency = 1;


//   %DCT2 = alloca [7 x i32], align 4, !MSB !129, !LSB !130, !extendFrom !129
ram_dual_port main_entry_DCT2 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_DCT2_address_a ),
	.wren_a( main_entry_DCT2_write_enable_a ),
	.data_a( main_entry_DCT2_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_DCT2_out_a ),
	.address_b( main_entry_DCT2_address_b ),
	.wren_b( main_entry_DCT2_write_enable_b ),
	.data_b( main_entry_DCT2_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_DCT2_out_b )
);
defparam main_entry_DCT2.width_a = 32;
defparam main_entry_DCT2.widthad_a = 3;
defparam main_entry_DCT2.width_be_a = 4;
defparam main_entry_DCT2.numwords_a = 7;
defparam main_entry_DCT2.width_b = 32;
defparam main_entry_DCT2.widthad_b = 3;
defparam main_entry_DCT2.width_be_b = 4;
defparam main_entry_DCT2.numwords_b = 7;
defparam main_entry_DCT2.latency = 1;


//   %DCT3 = alloca [7 x i32], align 4, !MSB !129, !LSB !130, !extendFrom !129
ram_dual_port main_entry_DCT3 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_DCT3_address_a ),
	.wren_a( main_entry_DCT3_write_enable_a ),
	.data_a( main_entry_DCT3_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_DCT3_out_a ),
	.address_b( main_entry_DCT3_address_b ),
	.wren_b( main_entry_DCT3_write_enable_b ),
	.data_b( main_entry_DCT3_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_DCT3_out_b )
);
defparam main_entry_DCT3.width_a = 32;
defparam main_entry_DCT3.widthad_a = 3;
defparam main_entry_DCT3.width_be_a = 4;
defparam main_entry_DCT3.numwords_a = 7;
defparam main_entry_DCT3.width_b = 32;
defparam main_entry_DCT3.widthad_b = 3;
defparam main_entry_DCT3.width_be_b = 4;
defparam main_entry_DCT3.numwords_b = 7;
defparam main_entry_DCT3.latency = 1;


//   %DCT4 = alloca [7 x i32], align 4, !MSB !129, !LSB !130, !extendFrom !129
ram_dual_port main_entry_DCT4 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_DCT4_address_a ),
	.wren_a( main_entry_DCT4_write_enable_a ),
	.data_a( main_entry_DCT4_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_DCT4_out_a ),
	.address_b( main_entry_DCT4_address_b ),
	.wren_b( main_entry_DCT4_write_enable_b ),
	.data_b( main_entry_DCT4_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_DCT4_out_b )
);
defparam main_entry_DCT4.width_a = 32;
defparam main_entry_DCT4.widthad_a = 3;
defparam main_entry_DCT4.width_be_a = 4;
defparam main_entry_DCT4.numwords_a = 7;
defparam main_entry_DCT4.width_b = 32;
defparam main_entry_DCT4.widthad_b = 3;
defparam main_entry_DCT4.width_be_b = 4;
defparam main_entry_DCT4.numwords_b = 7;
defparam main_entry_DCT4.latency = 1;


//   %DCT5 = alloca [7 x i32], align 4, !MSB !129, !LSB !130, !extendFrom !129
ram_dual_port main_entry_DCT5 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_DCT5_address_a ),
	.wren_a( main_entry_DCT5_write_enable_a ),
	.data_a( main_entry_DCT5_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_DCT5_out_a ),
	.address_b( main_entry_DCT5_address_b ),
	.wren_b( main_entry_DCT5_write_enable_b ),
	.data_b( main_entry_DCT5_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_DCT5_out_b )
);
defparam main_entry_DCT5.width_a = 32;
defparam main_entry_DCT5.widthad_a = 3;
defparam main_entry_DCT5.width_be_a = 4;
defparam main_entry_DCT5.numwords_a = 7;
defparam main_entry_DCT5.width_b = 32;
defparam main_entry_DCT5.widthad_b = 3;
defparam main_entry_DCT5.width_be_b = 4;
defparam main_entry_DCT5.numwords_b = 7;
defparam main_entry_DCT5.latency = 1;


//   %DCT6 = alloca [7 x i32], align 4, !MSB !129, !LSB !130, !extendFrom !129
ram_dual_port main_entry_DCT6 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_DCT6_address_a ),
	.wren_a( main_entry_DCT6_write_enable_a ),
	.data_a( main_entry_DCT6_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_DCT6_out_a ),
	.address_b( main_entry_DCT6_address_b ),
	.wren_b( main_entry_DCT6_write_enable_b ),
	.data_b( main_entry_DCT6_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_DCT6_out_b )
);
defparam main_entry_DCT6.width_a = 32;
defparam main_entry_DCT6.widthad_a = 3;
defparam main_entry_DCT6.width_be_a = 4;
defparam main_entry_DCT6.numwords_a = 7;
defparam main_entry_DCT6.width_b = 32;
defparam main_entry_DCT6.widthad_b = 3;
defparam main_entry_DCT6.width_be_b = 4;
defparam main_entry_DCT6.numwords_b = 7;
defparam main_entry_DCT6.latency = 1;


//   %DCT7 = alloca [7 x i32], align 4, !MSB !129, !LSB !130, !extendFrom !129
ram_dual_port main_entry_DCT7 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_DCT7_address_a ),
	.wren_a( main_entry_DCT7_write_enable_a ),
	.data_a( main_entry_DCT7_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_DCT7_out_a ),
	.address_b( main_entry_DCT7_address_b ),
	.wren_b( main_entry_DCT7_write_enable_b ),
	.data_b( main_entry_DCT7_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_DCT7_out_b )
);
defparam main_entry_DCT7.width_a = 32;
defparam main_entry_DCT7.widthad_a = 3;
defparam main_entry_DCT7.width_be_a = 4;
defparam main_entry_DCT7.numwords_a = 7;
defparam main_entry_DCT7.width_b = 32;
defparam main_entry_DCT7.widthad_b = 3;
defparam main_entry_DCT7.width_be_b = 4;
defparam main_entry_DCT7.numwords_b = 7;
defparam main_entry_DCT7.latency = 1;


//   %DCT8 = alloca [7 x i32], align 4, !MSB !129, !LSB !130, !extendFrom !129
ram_dual_port main_entry_DCT8 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_DCT8_address_a ),
	.wren_a( main_entry_DCT8_write_enable_a ),
	.data_a( main_entry_DCT8_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_DCT8_out_a ),
	.address_b( main_entry_DCT8_address_b ),
	.wren_b( main_entry_DCT8_write_enable_b ),
	.data_b( main_entry_DCT8_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_DCT8_out_b )
);
defparam main_entry_DCT8.width_a = 32;
defparam main_entry_DCT8.widthad_a = 3;
defparam main_entry_DCT8.width_be_a = 4;
defparam main_entry_DCT8.numwords_a = 7;
defparam main_entry_DCT8.width_b = 32;
defparam main_entry_DCT8.widthad_b = 3;
defparam main_entry_DCT8.width_be_b = 4;
defparam main_entry_DCT8.numwords_b = 7;
defparam main_entry_DCT8.latency = 1;

/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
	if (!fsm_stall) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("%d ", $signed(main_for_cond2_preheader_64_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_cond2_preheader_64_reg) === 1'bX) finish <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("%d ", $signed(main_for_cond2_preheader_63_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_cond2_preheader_63_reg) === 1'bX) finish <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("%d ", $signed(main_for_cond2_preheader_62_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_cond2_preheader_62_reg) === 1'bX) finish <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("%d ", $signed(main_for_cond2_preheader_61_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_cond2_preheader_61_reg) === 1'bX) finish <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("%d ", $signed(main_for_cond2_preheader_60_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_cond2_preheader_60_reg) === 1'bX) finish <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("%d ", $signed(main_for_cond2_preheader_59_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_cond2_preheader_59_reg) === 1'bX) finish <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("%d ", $signed(main_for_cond2_preheader_58_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_cond2_preheader_58_reg) === 1'bX) finish <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("%d ", $signed(main_for_cond2_preheader_57_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_cond2_preheader_57_reg) === 1'bX) finish <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_8)) begin
		$write("\n");
	end
end
/* synthesis translate_on */
always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  // synthesis parallel_case  
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_pipeline_wait_loop_2;
LEGUP_F_main_BB_for_cond2_preheader_8:
	if ((fsm_stall == 1'd0) && (main_for_cond2_preheader_exitcond1 == 1'd1))
		next_state = LEGUP_F_main_BB_for_end9_11;
	else if ((fsm_stall == 1'd0) && (main_for_cond2_preheader_exitcond1 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9;
LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10:
		next_state = LEGUP_F_main_BB_for_cond2_preheader_8;
LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9:
		next_state = LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10;
LEGUP_F_main_BB_for_cond2_preheader_preheader_3:
		next_state = LEGUP_F_main_BB_for_cond2_preheader_preheader_4;
LEGUP_F_main_BB_for_cond2_preheader_preheader_4:
		next_state = LEGUP_F_main_BB_for_cond2_preheader_preheader_5;
LEGUP_F_main_BB_for_cond2_preheader_preheader_5:
		next_state = LEGUP_F_main_BB_for_cond2_preheader_preheader_6;
LEGUP_F_main_BB_for_cond2_preheader_preheader_6:
		next_state = LEGUP_F_main_BB_for_cond2_preheader_preheader_7;
LEGUP_F_main_BB_for_cond2_preheader_preheader_7:
		next_state = LEGUP_F_main_BB_for_cond2_preheader_8;
LEGUP_F_main_BB_for_end9_11:
		next_state = LEGUP_0;
LEGUP_pipeline_wait_loop_2:
	if ((fsm_stall == 1'd0) && (loop_pipeline_finish == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond2_preheader_preheader_3;
	else if ((fsm_stall == 1'd0) && (loop_pipeline_finish == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond2_preheader_preheader_3;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
assign main_entry_0 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_0_reg <= main_entry_0;
	end
end
assign main_entry_1 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_1_reg <= main_entry_1;
	end
end
assign main_entry_2 = (1'd0 + (4 * 32'd1));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_2_reg <= main_entry_2;
	end
end
assign main_for_cond2_preheader_preheader_4 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_4_reg <= main_for_cond2_preheader_preheader_4;
	end
end
assign main_for_cond2_preheader_preheader_5 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_5_reg <= main_for_cond2_preheader_preheader_5;
	end
end
assign main_for_cond2_preheader_preheader_6 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_6_reg <= main_for_cond2_preheader_preheader_6;
	end
end
assign main_for_cond2_preheader_preheader_7 = (1'd0 + (4 * 32'd3));
assign main_for_cond2_preheader_preheader_8 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_8_reg <= main_for_cond2_preheader_preheader_8;
	end
end
assign main_for_cond2_preheader_preheader_9 = (1'd0 + (4 * 32'd1));
assign main_for_cond2_preheader_preheader_10 = (1'd0 + (4 * 32'd3));
assign main_for_cond2_preheader_preheader_11 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_11_reg <= main_for_cond2_preheader_preheader_11;
	end
end
assign main_for_cond2_preheader_preheader_12 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_12_reg <= main_for_cond2_preheader_preheader_12;
	end
end
assign main_for_cond2_preheader_preheader_13 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_13_reg <= main_for_cond2_preheader_preheader_13;
	end
end
assign main_for_cond2_preheader_preheader_14 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_14_reg <= main_for_cond2_preheader_preheader_14;
	end
end
assign main_for_cond2_preheader_preheader_15 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_15_reg <= main_for_cond2_preheader_preheader_15;
	end
end
assign main_for_cond2_preheader_preheader_16 = (1'd0 + (4 * 32'd3));
assign main_for_cond2_preheader_preheader_17 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_17_reg <= main_for_cond2_preheader_preheader_17;
	end
end
assign main_for_cond2_preheader_preheader_18 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_18_reg <= main_for_cond2_preheader_preheader_18;
	end
end
assign main_for_cond2_preheader_preheader_19 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_19_reg <= main_for_cond2_preheader_preheader_19;
	end
end
assign main_for_cond2_preheader_preheader_20 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_20_reg <= main_for_cond2_preheader_preheader_20;
	end
end
assign main_for_cond2_preheader_preheader_21 = (1'd0 + (4 * 32'd1));
assign main_for_cond2_preheader_preheader_22 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_22_reg <= main_for_cond2_preheader_preheader_22;
	end
end
assign main_for_cond2_preheader_preheader_23 = (1'd0 + (4 * 32'd3));
assign main_for_cond2_preheader_preheader_24 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_24_reg <= main_for_cond2_preheader_preheader_24;
	end
end
assign main_for_cond2_preheader_preheader_25 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_25_reg <= main_for_cond2_preheader_preheader_25;
	end
end
assign main_for_cond2_preheader_preheader_26 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_26_reg <= main_for_cond2_preheader_preheader_26;
	end
end
assign main_for_cond2_preheader_preheader_27 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_27_reg <= main_for_cond2_preheader_preheader_27;
	end
end
assign main_for_cond2_preheader_preheader_28 = (1'd0 + (4 * 32'd1));
assign main_for_cond2_preheader_preheader_29 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_29_reg <= main_for_cond2_preheader_preheader_29;
	end
end
assign main_for_cond2_preheader_preheader_30 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_30_reg <= main_for_cond2_preheader_preheader_30;
	end
end
assign main_for_cond2_preheader_preheader_31 = (1'd0 + (4 * 32'd1));
assign main_for_cond2_preheader_preheader_32 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_32_reg <= main_for_cond2_preheader_preheader_32;
	end
end
assign main_for_cond2_preheader_preheader_33 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_33_reg <= main_for_cond2_preheader_preheader_33;
	end
end
assign main_for_cond2_preheader_preheader_34 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_34_reg <= main_for_cond2_preheader_preheader_34;
	end
end
assign main_for_cond2_preheader_preheader_35 = (1'd0 + (4 * 32'd3));
assign main_for_cond2_preheader_preheader_36 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_36_reg <= main_for_cond2_preheader_preheader_36;
	end
end
assign main_for_cond2_preheader_preheader_37 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_37_reg <= main_for_cond2_preheader_preheader_37;
	end
end
assign main_for_cond2_preheader_preheader_38 = (1'd0 + (4 * 32'd1));
assign main_for_cond2_preheader_preheader_39 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_39_reg <= main_for_cond2_preheader_preheader_39;
	end
end
assign main_for_cond2_preheader_preheader_40 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_40_reg <= main_for_cond2_preheader_preheader_40;
	end
end
assign main_for_cond2_preheader_preheader_41 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_41_reg <= main_for_cond2_preheader_preheader_41;
	end
end
assign main_for_cond2_preheader_preheader_42 = (1'd0 + (4 * 32'd3));
assign main_for_cond2_preheader_preheader_43 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_43_reg <= main_for_cond2_preheader_preheader_43;
	end
end
assign main_for_cond2_preheader_preheader_44 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_44_reg <= main_for_cond2_preheader_preheader_44;
	end
end
assign main_for_cond2_preheader_preheader_45 = (1'd0 + (4 * 32'd1));
assign main_for_cond2_preheader_preheader_46 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_46_reg <= main_for_cond2_preheader_preheader_46;
	end
end
assign main_for_cond2_preheader_preheader_47 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_47_reg <= main_for_cond2_preheader_preheader_47;
	end
end
assign main_for_cond2_preheader_preheader_48 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_48_reg <= main_for_cond2_preheader_preheader_48;
	end
end
assign main_for_cond2_preheader_preheader_49 = (1'd0 + (4 * 32'd3));
assign main_for_cond2_preheader_preheader_50 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_50_reg <= main_for_cond2_preheader_preheader_50;
	end
end
assign main_for_cond2_preheader_preheader_51 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_51_reg <= main_for_cond2_preheader_preheader_51;
	end
end
assign main_for_cond2_preheader_preheader_52 = (1'd0 + (4 * 32'd1));
assign main_for_cond2_preheader_preheader_53 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_53_reg <= main_for_cond2_preheader_preheader_53;
	end
end
assign main_for_cond2_preheader_preheader_54 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_54_reg <= main_for_cond2_preheader_preheader_54;
	end
end
assign main_for_cond2_preheader_preheader_55 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_for_cond2_preheader_preheader_55_reg <= main_for_cond2_preheader_preheader_55;
	end
end
assign main_for_cond2_preheader_preheader_56 = (1'd0 + (4 * 32'd3));
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_57 = -32'd3;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_57 = main_for_cond2_preheader_for_cond2_preheader_crit__var15;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_57_reg <= main_for_cond2_preheader_57;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_57_reg <= main_for_cond2_preheader_57;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_58 = 32'd10;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_58 = main_for_cond2_preheader_for_cond2_preheader_crit__var14;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_58_reg <= main_for_cond2_preheader_58;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_58_reg <= main_for_cond2_preheader_58;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_59 = 32'd12;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_59 = main_for_cond2_preheader_for_cond2_preheader_crit__var13;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_59_reg <= main_for_cond2_preheader_59;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_59_reg <= main_for_cond2_preheader_59;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_60 = 32'd8;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_60 = main_for_cond2_preheader_for_cond2_preheader_crit__var12;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_60_reg <= main_for_cond2_preheader_60;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_60_reg <= main_for_cond2_preheader_60;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_61 = 32'd5;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_61 = main_for_cond2_preheader_for_cond2_preheader_crit__var11;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_61_reg <= main_for_cond2_preheader_61;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_61_reg <= main_for_cond2_preheader_61;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_62 = 32'd2;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_62 = main_for_cond2_preheader_for_cond2_preheader_crit__var10;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_62_reg <= main_for_cond2_preheader_62;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_62_reg <= main_for_cond2_preheader_62;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_63 = 32'd36;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_63 = main_for_cond2_preheader_for_cond2_preheader_crit__var9;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_63_reg <= main_for_cond2_preheader_63;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_63_reg <= main_for_cond2_preheader_63;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_64 = 32'd197;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_64 = main_for_cond2_preheader_for_cond2_preheader_crit__var8;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_64_reg <= main_for_cond2_preheader_64;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_64_reg <= main_for_cond2_preheader_64;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_65 = 32'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) */ begin
		main_for_cond2_preheader_65 = main_for_cond2_preheader_for_cond2_preheader_crit__var7_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_65_reg <= main_for_cond2_preheader_65;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_10) & (fsm_stall == 1'd0))) begin
		main_for_cond2_preheader_65_reg <= main_for_cond2_preheader_65;
	end
end
always @(*) begin
		main_for_cond2_preheader_exitcond1 = (main_for_cond2_preheader_65_reg == 32'd7);
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit_ = (1'd0 + (4 * {28'd0,main_for_cond2_preheader_65_reg}));
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var0 = (1'd0 + (4 * {28'd0,main_for_cond2_preheader_65_reg}));
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var1 = (1'd0 + (4 * {28'd0,main_for_cond2_preheader_65_reg}));
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var2 = (1'd0 + (4 * {28'd0,main_for_cond2_preheader_65_reg}));
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var3 = (1'd0 + (4 * {28'd0,main_for_cond2_preheader_65_reg}));
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var4 = (1'd0 + (4 * {28'd0,main_for_cond2_preheader_65_reg}));
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var5 = (1'd0 + (4 * {28'd0,main_for_cond2_preheader_65_reg}));
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var6 = (1'd0 + (4 * {28'd0,main_for_cond2_preheader_65_reg}));
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var7 = ({1'd0,main_for_cond2_preheader_65_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var7_reg <= main_for_cond2_preheader_for_cond2_preheader_crit__var7;
	end
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var8 = main_entry_DCT1_out_b;
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var9 = main_entry_DCT2_out_b;
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var10 = main_entry_DCT3_out_b;
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var11 = main_entry_DCT4_out_b;
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var12 = main_entry_DCT5_out_b;
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var13 = main_entry_DCT6_out_b;
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var14 = main_entry_DCT7_out_b;
end
always @(*) begin
		main_for_cond2_preheader_for_cond2_preheader_crit__var15 = main_entry_DCT8_out_b;
end
always @(*) begin
	main_entry_DCT1_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT1_address_a = (main_for_cond2_preheader_preheader_16 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT1_address_a = (main_for_cond2_preheader_preheader_8_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT1_address_a = (main_for_cond2_preheader_preheader_15_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT1_address_a = (main_for_cond2_preheader_preheader_4_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT1_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT1_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT1_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT1_in_a = 32'd27;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT1_in_a = -32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT1_in_a = -32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT1_in_a = -32'd24;
	end
end
always @(*) begin
	main_entry_DCT1_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT1_address_b = (main_for_cond2_preheader_preheader_31 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT1_address_b = (main_for_cond2_preheader_preheader_30_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT1_address_b = (main_for_cond2_preheader_preheader_29_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_entry_DCT1_address_b = (main_for_cond2_preheader_for_cond2_preheader_crit_ >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT1_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT1_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT1_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT1_in_b = 32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT1_in_b = 32'd20;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT1_in_b = -32'd12;
	end
end
always @(*) begin
	main_entry_DCT2_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT2_address_a = (main_for_cond2_preheader_preheader_35 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT2_address_a = (main_for_cond2_preheader_preheader_34_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT2_address_a = (main_for_cond2_preheader_preheader_33_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT2_address_a = (main_for_cond2_preheader_preheader_32_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT2_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT2_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT2_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT2_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT2_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT2_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT2_in_a = -32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT2_in_a = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT2_in_a = -32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT2_in_a = -32'd42;
	end
end
always @(*) begin
	main_entry_DCT2_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT2_address_b = (main_for_cond2_preheader_preheader_9 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT2_address_b = (main_for_cond2_preheader_preheader_17_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT2_address_b = (main_entry_0_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_entry_DCT2_address_b = (main_for_cond2_preheader_for_cond2_preheader_crit__var0 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT2_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT2_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT2_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT2_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT2_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT2_in_b = 32'd11;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT2_in_b = -32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT2_in_b = 32'd6;
	end
end
always @(*) begin
	main_entry_DCT3_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT3_address_a = (main_for_cond2_preheader_preheader_10 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT3_address_a = (main_for_cond2_preheader_preheader_19_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT3_address_a = (main_for_cond2_preheader_preheader_5_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT3_address_a = (main_for_cond2_preheader_preheader_18_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT3_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT3_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT3_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT3_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT3_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT3_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT3_in_a = -32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT3_in_a = -32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT3_in_a = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT3_in_a = -32'd22;
	end
end
always @(*) begin
	main_entry_DCT3_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT3_address_b = (main_for_cond2_preheader_preheader_38 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT3_address_b = (main_for_cond2_preheader_preheader_37_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT3_address_b = (main_for_cond2_preheader_preheader_36_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_entry_DCT3_address_b = (main_for_cond2_preheader_for_cond2_preheader_crit__var1 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT3_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT3_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT3_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT3_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT3_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT3_in_b = -32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT3_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT3_in_b = 32'd0;
	end
end
always @(*) begin
	main_entry_DCT4_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT4_address_a = (main_for_cond2_preheader_preheader_42 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT4_address_a = (main_for_cond2_preheader_preheader_41_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT4_address_a = (main_for_cond2_preheader_preheader_40_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT4_address_a = (main_for_cond2_preheader_preheader_39_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT4_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT4_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT4_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT4_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT4_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT4_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT4_in_a = -32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT4_in_a = -32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT4_in_a = -32'd13;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT4_in_a = -32'd12;
	end
end
always @(*) begin
	main_entry_DCT4_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT4_address_b = (main_for_cond2_preheader_preheader_21 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT4_address_b = (main_entry_1_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT4_address_b = (main_for_cond2_preheader_preheader_20_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_entry_DCT4_address_b = (main_for_cond2_preheader_for_cond2_preheader_crit__var2 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT4_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT4_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT4_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT4_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT4_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT4_in_b = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT4_in_b = -32'd7;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT4_in_b = -32'd6;
	end
end
always @(*) begin
	main_entry_DCT5_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT5_address_a = (main_for_cond2_preheader_preheader_23 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT5_address_a = (main_for_cond2_preheader_preheader_6_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT5_address_a = (main_for_cond2_preheader_preheader_22_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT5_address_a = (main_for_cond2_preheader_preheader_11_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT5_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT5_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT5_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT5_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT5_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT5_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT5_in_a = -32'd7;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT5_in_a = 32'd13;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT5_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT5_in_a = 32'd3;
	end
end
always @(*) begin
	main_entry_DCT5_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT5_address_b = (main_for_cond2_preheader_preheader_45 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT5_address_b = (main_for_cond2_preheader_preheader_44_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT5_address_b = (main_for_cond2_preheader_preheader_43_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_entry_DCT5_address_b = (main_for_cond2_preheader_for_cond2_preheader_crit__var3 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT5_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT5_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT5_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT5_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT5_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT5_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT5_in_b = -32'd14;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT5_in_b = 32'd14;
	end
end
always @(*) begin
	main_entry_DCT6_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT6_address_a = (main_for_cond2_preheader_preheader_49 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT6_address_a = (main_for_cond2_preheader_preheader_48_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT6_address_a = (main_for_cond2_preheader_preheader_47_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT6_address_a = (main_for_cond2_preheader_preheader_46_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT6_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT6_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT6_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT6_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT6_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT6_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT6_in_a = 32'd11;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT6_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT6_in_a = 32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT6_in_a = -32'd7;
	end
end
always @(*) begin
	main_entry_DCT6_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT6_address_b = (main_entry_2_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT6_address_b = (main_for_cond2_preheader_preheader_24_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT6_address_b = (main_for_cond2_preheader_preheader_12_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_entry_DCT6_address_b = (main_for_cond2_preheader_for_cond2_preheader_crit__var4 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT6_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT6_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT6_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT6_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT6_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT6_in_b = -32'd16;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT6_in_b = 32'd7;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT6_in_b = -32'd6;
	end
end
always @(*) begin
	main_entry_DCT7_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT7_address_a = (main_for_cond2_preheader_preheader_7 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT7_address_a = (main_for_cond2_preheader_preheader_26_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT7_address_a = (main_for_cond2_preheader_preheader_13_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT7_address_a = (main_for_cond2_preheader_preheader_25_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT7_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT7_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT7_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT7_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT7_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT7_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT7_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT7_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT7_in_a = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT7_in_a = -32'd2;
	end
end
always @(*) begin
	main_entry_DCT7_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT7_address_b = (main_for_cond2_preheader_preheader_52 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT7_address_b = (main_for_cond2_preheader_preheader_51_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT7_address_b = (main_for_cond2_preheader_preheader_50_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_entry_DCT7_address_b = (main_for_cond2_preheader_for_cond2_preheader_crit__var5 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT7_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT7_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT7_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT7_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT7_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT7_in_b = -32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT7_in_b = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT7_in_b = -32'd6;
	end
end
always @(*) begin
	main_entry_DCT8_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT8_address_a = (main_for_cond2_preheader_preheader_56 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT8_address_a = (main_for_cond2_preheader_preheader_55_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT8_address_a = (main_for_cond2_preheader_preheader_54_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT8_address_a = (main_for_cond2_preheader_preheader_53_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT8_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT8_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT8_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT8_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT8_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT8_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT8_in_a = -32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT8_in_a = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT8_in_a = -32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_6)) begin
		main_entry_DCT8_in_a = 32'd9;
	end
end
always @(*) begin
	main_entry_DCT8_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT8_address_b = (main_for_cond2_preheader_preheader_28 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT8_address_b = (main_for_cond2_preheader_preheader_14_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT8_address_b = (main_for_cond2_preheader_preheader_27_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_for_cond2_preheader_crit_edge_9)) begin
		main_entry_DCT8_address_b = (main_for_cond2_preheader_for_cond2_preheader_crit__var6 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_DCT8_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT8_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT8_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT8_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_DCT8_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_3)) begin
		main_entry_DCT8_in_b = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_4)) begin
		main_entry_DCT8_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond2_preheader_preheader_5)) begin
		main_entry_DCT8_in_b = -32'd3;
	end
end
always @(posedge clk) begin
	if (~(loop_state_stall_0)) begin
		loop_valid_bit_0 <= (loop_II_counter & loop_start);
	end
	if (reset) begin
		loop_valid_bit_0 <= 1'd0;
	end
end
assign loop_state_stall_0 = 1'd0;
always @(*) begin
	loop_state_enable_0 = (loop_valid_bit_0 & ~(loop_state_stall_0));
end
always @(posedge clk) begin
	loop_II_counter <= 1'd1;
end
always @(*) begin
	loop_start = (loop_activate_pipeline | ((loop_active & ~(loop_epilogue)) & ~((loop_state_enable_0 & loop_pipeline_exit_cond))));
	if (reset) begin
		loop_start = 1'd0;
	end
end
always @(*) begin
	loop_activate_pipeline = (((fsm_stall == 1'd0) & loop_begin_pipeline) & ~(loop_active));
end
always @(*) begin
	loop_pipeline_exit_cond = (loop_inductionVar_stage0 == 1583);
end
always @(posedge clk) begin
	if (reset) begin
		loop_inductionVar_stage0 <= 0;
	end
	if (loop_activate_pipeline) begin
		loop_inductionVar_stage0 <= 0;
	end
	if ((loop_II_counter & loop_state_enable_0)) begin
		loop_inductionVar_stage0 <= (loop_inductionVar_stage0 + 1'd1);
	end
end
always @(posedge clk) begin
	if (reset) begin
		loop_active <= 1'd0;
	end
	if (loop_activate_pipeline) begin
		loop_active <= 1'd1;
	end
	if ((loop_epilogue & loop_only_last_stage_enabled)) begin
		loop_active <= 1'd0;
	end
end
always @(*) begin
	loop_begin_pipeline = 1'd0;
	if (reset) begin
		loop_begin_pipeline = 1'd0;
	end
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		loop_begin_pipeline = 1'd1;
	end
end
always @(posedge clk) begin
	if (reset) begin
		loop_epilogue <= 1'd0;
	end
	if ((loop_state_enable_0 & loop_pipeline_exit_cond)) begin
		loop_epilogue <= 1'd1;
	end
	if ((loop_epilogue & loop_only_last_stage_enabled)) begin
		loop_epilogue <= 1'd0;
	end
end
always @(*) begin
	loop_pipeline_finish = ((loop_epilogue & loop_only_last_stage_enabled) | loop_pipeline_finish_reg);
end
always @(*) begin
	loop_only_last_stage_enabled = ~(loop_state_enable_0);
end
always @(posedge clk) begin
	loop_pipeline_finish_reg <= loop_pipeline_finish;
	if (reset) begin
		loop_pipeline_finish_reg <= 1'd0;
	end
	if (loop_activate_pipeline) begin
		loop_pipeline_finish_reg <= 1'd0;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end9_11)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end9_11)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
